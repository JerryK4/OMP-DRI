`timescale 1ns / 1ps

module finding_max(
    input wire clk,
    input wire rst_n,
    input wire start_search, 
    
    // Giao ti?p v?i Dot Product Engine
    input wire [47:0] dot_result,      
    input wire [5:0]  current_col_idx, 
    input wire        col_done,        
    input wire        all_done_in,     
    
    // Qu?n l� l?ch s? (Masking)
    input wire [4:0]   current_i,       
    input wire [111:0] lambda_history,  // 16 lambda x 7-bit
    
    // K?t qu? ??u ra
    output reg [5:0]  lambda,          
    output reg        finding_done     
);

    reg [47:0] max_val_reg;
    reg [5:0]  lambda_temp;
    reg        is_masked; 
    reg        first_valid_found; // C? b�o hi?u ?� t�m ???c c?t ??u ti�n kh�ng b? kh�a
    integer    k;

    // 1. T�nh gi� tr? tuy?t ??i (B?o to�n s? c� d?u Q20.26)
    wire [47:0] abs_val = dot_result[47] ? (~dot_result + 1'b1) : dot_result;

    // 2. Logic t�m Max v� Masking chu?n x�c
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            max_val_reg <= 48'd0;
            lambda_temp <= 6'd0;
            lambda      <= 6'd0;
            finding_done <= 1'b0;
            first_valid_found <= 1'b0;
        end else begin
            if (start_search) begin
                // Reset tr?ng th�i cho ??t t�m ki?m m?i trong v�ng l?p OMP hi?n t?i
                max_val_reg <= 48'd0;
                lambda_temp <= 6'd0;
                finding_done <= 1'b0;
                first_valid_found <= 1'b0;
            end 
            else if (col_done) begin
                // --- B??C 1: KI?M TRA MASKING ---
                is_masked = 0; // Blocking assignment ?? c� k?t qu? ngay cho if ph�a d??i
                for (k = 0; k < 16; k = k + 1) begin
                    if (k < current_i) begin
                        // Ki?m tra: Tr�ng index V� � nh? history ?� ph?i h?p l? (bit[6] == 0)
                        if (current_col_idx == lambda_history[k*7 +: 6] && lambda_history[k*7 + 6] == 1'b0)
                            is_masked = 1;
                    end
                end

                // --- B??C 2: SO S�NH T�M MAX ---
                if (!is_masked) begin
                    // N?u ?�y l� c?t h?p l? (kh�ng b? mask) ??u ti�n t�m th?y
                    if (!first_valid_found) begin
                        max_val_reg <= abs_val;
                        lambda_temp <= current_col_idx;
                        first_valid_found <= 1'b1;
                    end
                    // Ho?c n?u t�m th?y c?t c� ?? t??ng quan th?c s? l?n h?n c?t Max c?
                    else if (abs_val > max_val_reg) begin
                        max_val_reg <= abs_val;
                        lambda_temp <= current_col_idx;
                    end
                end
            end 
            
            // --- B??C 3: CH?T K?T QU? ---
            if (all_done_in) begin
                lambda <= lambda_temp;
                finding_done <= 1'b1;
            end else begin
                finding_done <= 1'b0;
            end 
        end
    end

endmodule